PO4A-HEADER: mode=after; position=F�RFATTARE; beginboundary=\.SH
.SH �VERS�TTARE
Denna manualsida har �versatts av Daniel Nylander <po@danielnylander.se> 
den 31 oktober 2005.

Om du hittar n�gra felaktigheter i �vers�ttningen, v�nligen skicka ett 
e-postmeddelande till �versättaren eller till e-postlistan
.nh
<\fIdebian\-l10n\-swedish@lists.debian.org\fR> eller <\fItp-sv@listor.tp-sv.se\fR>
.hy

